module Small_FV_MEMCntl(

    
);


endmodule


